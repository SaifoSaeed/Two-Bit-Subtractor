module XOR_G(
    x,
    y,
    z
);

input wire x, y;
output wire z;

assign z = x ^ y;
    
endmodule